*** SPICE deck for cell carry-out-2x{sch} from library carry-out-2x
*** Created on Tue Sep 26, 2023 22:59:56
*** Last revised on Fri Oct 27, 2023 12:47:49
*** Written on Fri Oct 27, 2023 13:52:42 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: carry-out-2x{sch}
Mnmos@0 net@0 A gnd gnd nmos L=0.022U W=0.088U
Mnmos@1 net@0 A gnd gnd nmos L=0.022U W=0.088U
Mnmos@3 net@0 B gnd gnd nmos L=0.022U W=0.088U
Mnmos@4 net@0 B gnd gnd nmos L=0.022U W=0.088U
Mnmos@6 Y C net@0 gnd nmos L=0.022U W=0.088U
Mnmos@7 Y C net@0 gnd nmos L=0.022U W=0.088U
Mnmos@9 Y A net@41 gnd nmos L=0.022U W=0.088U
Mnmos@10 net@41 B gnd gnd nmos L=0.022U W=0.088U
Mpmos@0 vdd A net@53 vdd pmos L=0.022U W=0.176U
Mpmos@1 vdd A net@53 vdd pmos L=0.022U W=0.176U
Mpmos@3 vdd B net@53 vdd pmos L=0.022U W=0.176U
Mpmos@4 vdd B net@53 vdd pmos L=0.022U W=0.176U
Mpmos@6 net@53 C Y vdd pmos L=0.022U W=0.176U
Mpmos@7 net@53 C Y vdd pmos L=0.022U W=0.176U
Mpmos@9 vdd B net@40 vdd pmos L=0.022U W=0.176U
Mpmos@10 net@40 A Y vdd pmos L=0.022U W=0.176U

* Spice Code nodes in cell cell 'carry-out-2x{sch}'
.include "C:\Users\ganga\OneDrive\Desktop\DIC\22nm_HP.pm"
.param vdd = 0.8
v1 vdd gnd DC {vdd}
v2 A gnd PULSE(0 {vdd} 100p 100p 100p 700p 2n)
v3 B gnd PULSE(0 {vdd} 100p 100p 100p 350p 1n)
v4 C gnd PULSE(0 {vdd} 100p 100p 100p 175p 1n)
.meas tran delay_a_to_y
+trig v(a) val = (vdd/2) cross = 2
+targ v(y) val = (vdd/2) cross = 2
.tran 0 2n
.END
.END
